temporayr file

new feature added