temporayr file

new feature added (switch)
want to go prev version
