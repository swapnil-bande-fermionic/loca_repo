temporayr file

new feature added (switch)