temporayr file

new feature added (stch)
