temporayr file