temporayr file

new feature added (button)